* AVE SPICE Model: L-Alanine
* Backbone topology mapped to L/C tensors

* --- The Amino Source (NH3+) ---
V_amino in 0 SIN(0 1V 100GHz)
L_nh3 in n_amino 140.07pH
C_nc n_amino n_alpha 170.64846416382252fF

* --- The Alpha Carbon (C-alpha) ---
L_alpha n_alpha n_alpha_out 120.10999999999999pH

* --- R-Group Filter Stub (L-Alanine) ---
C_rgroup_bond n_alpha n_r_carbon 144.0922190201729fF
L_r_carbon n_r_carbon n_r_h_split 120.10999999999999pH
C_ch1 n_r_h_split n_rh1 121.06537530266344fF
L_rh1 n_rh1 0 10.08pH
C_ch2 n_r_h_split n_rh2 121.06537530266344fF
L_rh2 n_rh2 0 10.08pH
C_ch3 n_r_h_split n_rh3 121.06537530266344fF
L_rh3 n_rh3 0 10.08pH

C_cc n_alpha_out n_carboxyl_c 144.0922190201729fF

* --- The Carboxyl Sink (COO-) ---
L_carboxyl_c n_carboxyl_c n_carboxyl_split 120.10999999999999pH
C_co_double n_carboxyl_split n_o_double 62.57822277847309fF
L_o_double n_o_double 0 159.99pH
C_co_single n_carboxyl_split out 139.66480446927375fF
L_o_single out n_term 159.99pH
R_load n_term 0 376.73Ohm

* --- AC Simulation Directives ---
.ac dec 100 1G 1000G
.end
