* AVE SPICE Model: L-Alanine
* Backbone topology mapped to L/C tensors

* --- The Amino Source (NH3+) ---
V_amino in 0 SIN(0 1V 30THz)
L_nh3 in n_amino 1.3511297647809685e-13pH
C_nc n_amino n_alpha 3.9499212740708347e-16fF

* --- The Alpha Carbon (C-alpha) ---
L_alpha n_alpha n_alpha_out 1.1585894083442053e-13pH

* --- R-Group Filter Stub (L-Alanine) ---
C_rgroup_bond n_alpha n_r_carbon 4.576118317492612e-16fF
L_r_carbon n_r_carbon n_r_h_split 1.1585894083442053e-13pH
C_ch1 n_r_h_split n_rh1 3.6465177285491996e-16fF
L_rh1 n_rh1 0 9.72290214763884e-15pH
C_ch2 n_r_h_split n_rh2 3.6465177285491996e-16fF
L_rh2 n_rh2 0 9.72290214763884e-15pH
C_ch3 n_r_h_split n_rh3 3.6465177285491996e-16fF
L_rh3 n_rh3 0 9.72290214763884e-15pH

C_cc n_alpha_out n_carboxyl_c 4.576118317492612e-16fF

* --- The Carboxyl Sink (COO-) ---
L_carboxyl_c n_carboxyl_c n_carboxyl_split 1.1585894083442053e-13pH
C_co_double n_carboxyl_split n_o_double 1.2854565915673514e-16fF
L_o_double n_o_double 0 1.543351792973122e-13pH
C_co_single n_carboxyl_split out 3.5540363769155313e-16fF
L_o_single out n_term 1.543351792973122e-13pH
R_load n_term 0 376.7303Ohm

* --- AC Simulation Directives ---
.ac dec 100 1G 1000G
.end
