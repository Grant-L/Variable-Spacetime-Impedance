* Applied Vacuum Engineering - PONDER-01 Testbench
* Asymmetric AC Geometry: Carbon-12 Emitter vs Flat Collector



* -----------------------------------------------------------------
* NUCLEON (Baseline 6^3_2 Topological Defect)
* -----------------------------------------------------------------
.SUBCKT NUCLEON IN OUT
L_CORE IN OUT 1uH
C_CORE IN OUT 1pF
.ENDS NUCLEON



* -----------------------------------------------------------------
* MACROSCOPIC TOPOLOGY
* -----------------------------------------------------------------
V_VHF NODE_E 0 AC 1 SINE(0 30k 100MEG)

X_EMIT_1 NODE_E 0 NUCLEON
X_EMIT_2 NODE_E 0 NUCLEON
X_EMIT_3 NODE_E 0 NUCLEON
X_EMIT_4 NODE_E 0 NUCLEON
X_EMIT_5 NODE_E 0 NUCLEON
X_EMIT_6 NODE_E 0 NUCLEON
X_EMIT_7 NODE_E 0 NUCLEON
X_EMIT_8 NODE_E 0 NUCLEON
X_EMIT_9 NODE_E 0 NUCLEON
X_EMIT_10 NODE_E 0 NUCLEON
X_EMIT_11 NODE_E 0 NUCLEON
X_EMIT_12 NODE_E 0 NUCLEON
X_COLL_1 0 0 NUCLEON
X_COLL_2 0 0 NUCLEON
X_COLL_3 0 0 NUCLEON
X_COLL_4 0 0 NUCLEON
X_COLL_5 0 0 NUCLEON
X_COLL_6 0 0 NUCLEON
X_COLL_7 0 0 NUCLEON
X_COLL_8 0 0 NUCLEON
X_COLL_9 0 0 NUCLEON


* -----------------------------------------------------------------
* SPATIAL MUTUAL INDUCTANCE (K-FACTORS)
* -----------------------------------------------------------------
K_1 X_EMIT_1.L_CORE X_EMIT_2.L_CORE 0.207973
K_2 X_EMIT_1.L_CORE X_EMIT_3.L_CORE 0.207973
K_3 X_EMIT_1.L_CORE X_EMIT_4.L_CORE 0.207973
K_4 X_EMIT_1.L_CORE X_EMIT_5.L_CORE 0.006683
K_5 X_EMIT_1.L_CORE X_EMIT_6.L_CORE 0.006625
K_6 X_EMIT_1.L_CORE X_EMIT_7.L_CORE 0.006552
K_7 X_EMIT_1.L_CORE X_EMIT_8.L_CORE 0.006756
K_8 X_EMIT_1.L_CORE X_EMIT_9.L_CORE 0.006683
K_9 X_EMIT_1.L_CORE X_EMIT_10.L_CORE 0.006481
K_10 X_EMIT_1.L_CORE X_EMIT_11.L_CORE 0.006552
K_11 X_EMIT_1.L_CORE X_EMIT_12.L_CORE 0.006605
K_12 X_EMIT_2.L_CORE X_EMIT_3.L_CORE 0.207973
K_13 X_EMIT_2.L_CORE X_EMIT_4.L_CORE 0.207973
K_14 X_EMIT_2.L_CORE X_EMIT_5.L_CORE 0.006736
K_15 X_EMIT_2.L_CORE X_EMIT_6.L_CORE 0.006683
K_16 X_EMIT_2.L_CORE X_EMIT_7.L_CORE 0.006605
K_17 X_EMIT_2.L_CORE X_EMIT_8.L_CORE 0.006815
K_18 X_EMIT_2.L_CORE X_EMIT_9.L_CORE 0.006897
K_19 X_EMIT_2.L_CORE X_EMIT_10.L_CORE 0.006683
K_20 X_EMIT_2.L_CORE X_EMIT_11.L_CORE 0.006756
K_21 X_EMIT_2.L_CORE X_EMIT_12.L_CORE 0.006815
K_22 X_EMIT_3.L_CORE X_EMIT_4.L_CORE 0.207973
K_23 X_EMIT_3.L_CORE X_EMIT_5.L_CORE 0.006815
K_24 X_EMIT_3.L_CORE X_EMIT_6.L_CORE 0.006756
K_25 X_EMIT_3.L_CORE X_EMIT_7.L_CORE 0.006683
K_26 X_EMIT_3.L_CORE X_EMIT_8.L_CORE 0.006897
K_27 X_EMIT_3.L_CORE X_EMIT_9.L_CORE 0.006815
K_28 X_EMIT_3.L_CORE X_EMIT_10.L_CORE 0.006605
K_29 X_EMIT_3.L_CORE X_EMIT_11.L_CORE 0.006683
K_30 X_EMIT_3.L_CORE X_EMIT_12.L_CORE 0.006736
K_31 X_EMIT_4.L_CORE X_EMIT_5.L_CORE 0.006605
K_32 X_EMIT_4.L_CORE X_EMIT_6.L_CORE 0.006552
K_33 X_EMIT_4.L_CORE X_EMIT_7.L_CORE 0.006481
K_34 X_EMIT_4.L_CORE X_EMIT_8.L_CORE 0.006683
K_35 X_EMIT_4.L_CORE X_EMIT_9.L_CORE 0.006756
K_36 X_EMIT_4.L_CORE X_EMIT_10.L_CORE 0.006552
K_37 X_EMIT_4.L_CORE X_EMIT_11.L_CORE 0.006625
K_38 X_EMIT_4.L_CORE X_EMIT_12.L_CORE 0.006683
K_39 X_EMIT_5.L_CORE X_EMIT_6.L_CORE 0.207973
K_40 X_EMIT_5.L_CORE X_EMIT_7.L_CORE 0.207973
K_41 X_EMIT_5.L_CORE X_EMIT_8.L_CORE 0.207973
K_42 X_EMIT_5.L_CORE X_EMIT_9.L_CORE 0.006683
K_43 X_EMIT_5.L_CORE X_EMIT_10.L_CORE 0.006533
K_44 X_EMIT_5.L_CORE X_EMIT_11.L_CORE 0.006679
K_45 X_EMIT_5.L_CORE X_EMIT_12.L_CORE 0.006533
K_46 X_EMIT_6.L_CORE X_EMIT_7.L_CORE 0.207973
K_47 X_EMIT_6.L_CORE X_EMIT_8.L_CORE 0.207973
K_48 X_EMIT_6.L_CORE X_EMIT_9.L_CORE 0.006836
K_49 X_EMIT_6.L_CORE X_EMIT_10.L_CORE 0.006683
K_50 X_EMIT_6.L_CORE X_EMIT_11.L_CORE 0.006836
K_51 X_EMIT_6.L_CORE X_EMIT_12.L_CORE 0.006679
K_52 X_EMIT_7.L_CORE X_EMIT_8.L_CORE 0.207973
K_53 X_EMIT_7.L_CORE X_EMIT_9.L_CORE 0.006679
K_54 X_EMIT_7.L_CORE X_EMIT_10.L_CORE 0.006533
K_55 X_EMIT_7.L_CORE X_EMIT_11.L_CORE 0.006683
K_56 X_EMIT_7.L_CORE X_EMIT_12.L_CORE 0.006533
K_57 X_EMIT_8.L_CORE X_EMIT_9.L_CORE 0.006836
K_58 X_EMIT_8.L_CORE X_EMIT_10.L_CORE 0.006679
K_59 X_EMIT_8.L_CORE X_EMIT_11.L_CORE 0.006836
K_60 X_EMIT_8.L_CORE X_EMIT_12.L_CORE 0.006683
K_61 X_EMIT_9.L_CORE X_EMIT_10.L_CORE 0.207973
K_62 X_EMIT_9.L_CORE X_EMIT_11.L_CORE 0.207973
K_63 X_EMIT_9.L_CORE X_EMIT_12.L_CORE 0.207973
K_64 X_EMIT_10.L_CORE X_EMIT_11.L_CORE 0.207973
K_65 X_EMIT_10.L_CORE X_EMIT_12.L_CORE 0.207973
K_66 X_EMIT_11.L_CORE X_EMIT_12.L_CORE 0.207973
K_67 X_COLL_1.L_CORE X_COLL_2.L_CORE 0.117647
K_68 X_COLL_1.L_CORE X_COLL_3.L_CORE 0.058824
K_69 X_COLL_1.L_CORE X_COLL_4.L_CORE 0.117647
K_70 X_COLL_1.L_CORE X_COLL_5.L_CORE 0.083189
K_71 X_COLL_1.L_CORE X_COLL_6.L_CORE 0.052613
K_72 X_COLL_1.L_CORE X_COLL_7.L_CORE 0.058824
K_73 X_COLL_1.L_CORE X_COLL_8.L_CORE 0.052613
K_74 X_COLL_1.L_CORE X_COLL_9.L_CORE 0.041595
K_75 X_COLL_2.L_CORE X_COLL_3.L_CORE 0.117647
K_76 X_COLL_2.L_CORE X_COLL_4.L_CORE 0.083189
K_77 X_COLL_2.L_CORE X_COLL_5.L_CORE 0.117647
K_78 X_COLL_2.L_CORE X_COLL_6.L_CORE 0.083189
K_79 X_COLL_2.L_CORE X_COLL_7.L_CORE 0.052613
K_80 X_COLL_2.L_CORE X_COLL_8.L_CORE 0.058824
K_81 X_COLL_2.L_CORE X_COLL_9.L_CORE 0.052613
K_82 X_COLL_3.L_CORE X_COLL_4.L_CORE 0.052613
K_83 X_COLL_3.L_CORE X_COLL_5.L_CORE 0.083189
K_84 X_COLL_3.L_CORE X_COLL_6.L_CORE 0.117647
K_85 X_COLL_3.L_CORE X_COLL_7.L_CORE 0.041595
K_86 X_COLL_3.L_CORE X_COLL_8.L_CORE 0.052613
K_87 X_COLL_3.L_CORE X_COLL_9.L_CORE 0.058824
K_88 X_COLL_4.L_CORE X_COLL_5.L_CORE 0.117647
K_89 X_COLL_4.L_CORE X_COLL_6.L_CORE 0.058824
K_90 X_COLL_4.L_CORE X_COLL_7.L_CORE 0.117647
K_91 X_COLL_4.L_CORE X_COLL_8.L_CORE 0.083189
K_92 X_COLL_4.L_CORE X_COLL_9.L_CORE 0.052613
K_93 X_COLL_5.L_CORE X_COLL_6.L_CORE 0.117647
K_94 X_COLL_5.L_CORE X_COLL_7.L_CORE 0.083189
K_95 X_COLL_5.L_CORE X_COLL_8.L_CORE 0.117647
K_96 X_COLL_5.L_CORE X_COLL_9.L_CORE 0.083189
K_97 X_COLL_6.L_CORE X_COLL_7.L_CORE 0.052613
K_98 X_COLL_6.L_CORE X_COLL_8.L_CORE 0.083189
K_99 X_COLL_6.L_CORE X_COLL_9.L_CORE 0.117647
K_100 X_COLL_7.L_CORE X_COLL_8.L_CORE 0.117647
K_101 X_COLL_7.L_CORE X_COLL_9.L_CORE 0.058824
K_102 X_COLL_8.L_CORE X_COLL_9.L_CORE 0.117647
* -- Rectification Gradient (Gap Trans-Admittance) --
K_103 X_EMIT_1.L_CORE X_COLL_1.L_CORE 0.007681
K_104 X_EMIT_1.L_CORE X_COLL_2.L_CORE 0.007704
K_105 X_EMIT_1.L_CORE X_COLL_3.L_CORE 0.007694
K_106 X_EMIT_1.L_CORE X_COLL_4.L_CORE 0.008063
K_107 X_EMIT_1.L_CORE X_COLL_5.L_CORE 0.008090
K_108 X_EMIT_1.L_CORE X_COLL_6.L_CORE 0.008078
K_109 X_EMIT_1.L_CORE X_COLL_7.L_CORE 0.008465
K_110 X_EMIT_1.L_CORE X_COLL_8.L_CORE 0.008496
K_111 X_EMIT_1.L_CORE X_COLL_9.L_CORE 0.008482
K_112 X_EMIT_2.L_CORE X_COLL_1.L_CORE 0.007845
K_113 X_EMIT_2.L_CORE X_COLL_2.L_CORE 0.007856
K_114 X_EMIT_2.L_CORE X_COLL_3.L_CORE 0.007831
K_115 X_EMIT_2.L_CORE X_COLL_4.L_CORE 0.008238
K_116 X_EMIT_2.L_CORE X_COLL_5.L_CORE 0.008250
K_117 X_EMIT_2.L_CORE X_COLL_6.L_CORE 0.008222
K_118 X_EMIT_2.L_CORE X_COLL_7.L_CORE 0.008649
K_119 X_EMIT_2.L_CORE X_COLL_8.L_CORE 0.008663
K_120 X_EMIT_2.L_CORE X_COLL_9.L_CORE 0.008630
K_121 X_EMIT_3.L_CORE X_COLL_1.L_CORE 0.007974
K_122 X_EMIT_3.L_CORE X_COLL_2.L_CORE 0.008000
K_123 X_EMIT_3.L_CORE X_COLL_3.L_CORE 0.007988
K_124 X_EMIT_3.L_CORE X_COLL_4.L_CORE 0.008387
K_125 X_EMIT_3.L_CORE X_COLL_5.L_CORE 0.008417
K_126 X_EMIT_3.L_CORE X_COLL_6.L_CORE 0.008404
K_127 X_EMIT_3.L_CORE X_COLL_7.L_CORE 0.008822
K_128 X_EMIT_3.L_CORE X_COLL_8.L_CORE 0.008857
K_129 X_EMIT_3.L_CORE X_COLL_9.L_CORE 0.008842
K_130 X_EMIT_4.L_CORE X_COLL_1.L_CORE 0.007829
K_131 X_EMIT_4.L_CORE X_COLL_2.L_CORE 0.007839
K_132 X_EMIT_4.L_CORE X_COLL_3.L_CORE 0.007815
K_133 X_EMIT_4.L_CORE X_COLL_4.L_CORE 0.008235
K_134 X_EMIT_4.L_CORE X_COLL_5.L_CORE 0.008247
K_135 X_EMIT_4.L_CORE X_COLL_6.L_CORE 0.008219
K_136 X_EMIT_4.L_CORE X_COLL_7.L_CORE 0.008665
K_137 X_EMIT_4.L_CORE X_COLL_8.L_CORE 0.008679
K_138 X_EMIT_4.L_CORE X_COLL_9.L_CORE 0.008646
K_139 X_EMIT_5.L_CORE X_COLL_1.L_CORE 0.007947
K_140 X_EMIT_5.L_CORE X_COLL_2.L_CORE 0.008316
K_141 X_EMIT_5.L_CORE X_COLL_3.L_CORE 0.008693
K_142 X_EMIT_5.L_CORE X_COLL_4.L_CORE 0.007793
K_143 X_EMIT_5.L_CORE X_COLL_5.L_CORE 0.008139
K_144 X_EMIT_5.L_CORE X_COLL_6.L_CORE 0.008492
K_145 X_EMIT_5.L_CORE X_COLL_7.L_CORE 0.007615
K_146 X_EMIT_5.L_CORE X_COLL_8.L_CORE 0.007938
K_147 X_EMIT_5.L_CORE X_COLL_9.L_CORE 0.008264
K_148 X_EMIT_6.L_CORE X_COLL_1.L_CORE 0.008031
K_149 X_EMIT_6.L_CORE X_COLL_2.L_CORE 0.008395
K_150 X_EMIT_6.L_CORE X_COLL_3.L_CORE 0.008765
K_151 X_EMIT_6.L_CORE X_COLL_4.L_CORE 0.007858
K_152 X_EMIT_6.L_CORE X_COLL_5.L_CORE 0.008198
K_153 X_EMIT_6.L_CORE X_COLL_6.L_CORE 0.008541
K_154 X_EMIT_6.L_CORE X_COLL_7.L_CORE 0.007663
K_155 X_EMIT_6.L_CORE X_COLL_8.L_CORE 0.007977
K_156 X_EMIT_6.L_CORE X_COLL_9.L_CORE 0.008292
K_157 X_EMIT_7.L_CORE X_COLL_1.L_CORE 0.008034
K_158 X_EMIT_7.L_CORE X_COLL_2.L_CORE 0.008416
K_159 X_EMIT_7.L_CORE X_COLL_3.L_CORE 0.008808
K_160 X_EMIT_7.L_CORE X_COLL_4.L_CORE 0.007861
K_161 X_EMIT_7.L_CORE X_COLL_5.L_CORE 0.008217
K_162 X_EMIT_7.L_CORE X_COLL_6.L_CORE 0.008581
K_163 X_EMIT_7.L_CORE X_COLL_7.L_CORE 0.007666
K_164 X_EMIT_7.L_CORE X_COLL_8.L_CORE 0.007995
K_165 X_EMIT_7.L_CORE X_COLL_9.L_CORE 0.008329
K_166 X_EMIT_8.L_CORE X_COLL_1.L_CORE 0.008251
K_167 X_EMIT_8.L_CORE X_COLL_2.L_CORE 0.008647
K_168 X_EMIT_8.L_CORE X_COLL_3.L_CORE 0.009052
K_169 X_EMIT_8.L_CORE X_COLL_4.L_CORE 0.008079
K_170 X_EMIT_8.L_CORE X_COLL_5.L_CORE 0.008449
K_171 X_EMIT_8.L_CORE X_COLL_6.L_CORE 0.008826
K_172 X_EMIT_8.L_CORE X_COLL_7.L_CORE 0.007881
K_173 X_EMIT_8.L_CORE X_COLL_8.L_CORE 0.008224
K_174 X_EMIT_8.L_CORE X_COLL_9.L_CORE 0.008570
K_175 X_EMIT_9.L_CORE X_COLL_1.L_CORE 0.008845
K_176 X_EMIT_9.L_CORE X_COLL_2.L_CORE 0.008466
K_177 X_EMIT_9.L_CORE X_COLL_3.L_CORE 0.008093
K_178 X_EMIT_9.L_CORE X_COLL_4.L_CORE 0.008634
K_179 X_EMIT_9.L_CORE X_COLL_5.L_CORE 0.008280
K_180 X_EMIT_9.L_CORE X_COLL_6.L_CORE 0.007930
K_181 X_EMIT_9.L_CORE X_COLL_7.L_CORE 0.008394
K_182 X_EMIT_9.L_CORE X_COLL_8.L_CORE 0.008068
K_183 X_EMIT_9.L_CORE X_COLL_9.L_CORE 0.007743
K_184 X_EMIT_10.L_CORE X_COLL_1.L_CORE 0.008617
K_185 X_EMIT_10.L_CORE X_COLL_2.L_CORE 0.008249
K_186 X_EMIT_10.L_CORE X_COLL_3.L_CORE 0.007888
K_187 X_EMIT_10.L_CORE X_COLL_4.L_CORE 0.008404
K_188 X_EMIT_10.L_CORE X_COLL_5.L_CORE 0.008061
K_189 X_EMIT_10.L_CORE X_COLL_6.L_CORE 0.007724
K_190 X_EMIT_10.L_CORE X_COLL_7.L_CORE 0.008166
K_191 X_EMIT_10.L_CORE X_COLL_8.L_CORE 0.007851
K_192 X_EMIT_10.L_CORE X_COLL_9.L_CORE 0.007539
K_193 X_EMIT_11.L_CORE X_COLL_1.L_CORE 0.008966
K_194 X_EMIT_11.L_CORE X_COLL_2.L_CORE 0.008572
K_195 X_EMIT_11.L_CORE X_COLL_3.L_CORE 0.008185
K_196 X_EMIT_11.L_CORE X_COLL_4.L_CORE 0.008727
K_197 X_EMIT_11.L_CORE X_COLL_5.L_CORE 0.008362
K_198 X_EMIT_11.L_CORE X_COLL_6.L_CORE 0.008002
K_199 X_EMIT_11.L_CORE X_COLL_7.L_CORE 0.008462
K_200 X_EMIT_11.L_CORE X_COLL_8.L_CORE 0.008128
K_201 X_EMIT_11.L_CORE X_COLL_9.L_CORE 0.007796
K_202 X_EMIT_12.L_CORE X_COLL_1.L_CORE 0.008890
K_203 X_EMIT_12.L_CORE X_COLL_2.L_CORE 0.008487
K_204 X_EMIT_12.L_CORE X_COLL_3.L_CORE 0.008096
K_205 X_EMIT_12.L_CORE X_COLL_4.L_CORE 0.008675
K_206 X_EMIT_12.L_CORE X_COLL_5.L_CORE 0.008300
K_207 X_EMIT_12.L_CORE X_COLL_6.L_CORE 0.007933
K_208 X_EMIT_12.L_CORE X_COLL_7.L_CORE 0.008432
K_209 X_EMIT_12.L_CORE X_COLL_8.L_CORE 0.008086
K_210 X_EMIT_12.L_CORE X_COLL_9.L_CORE 0.007746


* -----------------------------------------------------------------
* SIMULATION DIRECTIVES
* -----------------------------------------------------------------
.TRAN 0.1n 50n
* Monitor the inductive momentum coupling across the gap
.PROBE V(NODE_E)

.END
