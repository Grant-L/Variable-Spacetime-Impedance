* Applied Vacuum Engineering - PONDER-01 Testbench
* Asymmetric AC Geometry: Helium-4 Emitter vs Flat Collector



* -----------------------------------------------------------------
* NUCLEON (Baseline 6^3_2 Topological Defect)
* -----------------------------------------------------------------
.SUBCKT NUCLEON IN OUT
L_CORE IN OUT 1uH
C_CORE IN OUT 1pF
.ENDS NUCLEON



* -----------------------------------------------------------------
* MACROSCOPIC TOPOLOGY
* -----------------------------------------------------------------
V_VHF NODE_E 0 AC 1 SINE(0 30k 100MEG)

X_EMIT_1 NODE_E 0 NUCLEON
X_EMIT_2 NODE_E 0 NUCLEON
X_EMIT_3 NODE_E 0 NUCLEON
X_EMIT_4 NODE_E 0 NUCLEON
X_COLL_1 0 0 NUCLEON
X_COLL_2 0 0 NUCLEON
X_COLL_3 0 0 NUCLEON
X_COLL_4 0 0 NUCLEON
X_COLL_5 0 0 NUCLEON
X_COLL_6 0 0 NUCLEON
X_COLL_7 0 0 NUCLEON
X_COLL_8 0 0 NUCLEON
X_COLL_9 0 0 NUCLEON


* -----------------------------------------------------------------
* SPATIAL MUTUAL INDUCTANCE (K-FACTORS)
* -----------------------------------------------------------------
K_1 X_EMIT_1.L_CORE X_EMIT_2.L_CORE 0.207973
K_2 X_EMIT_1.L_CORE X_EMIT_3.L_CORE 0.207973
K_3 X_EMIT_1.L_CORE X_EMIT_4.L_CORE 0.207973
K_4 X_EMIT_2.L_CORE X_EMIT_3.L_CORE 0.207973
K_5 X_EMIT_2.L_CORE X_EMIT_4.L_CORE 0.207973
K_6 X_EMIT_3.L_CORE X_EMIT_4.L_CORE 0.207973
K_7 X_COLL_1.L_CORE X_COLL_2.L_CORE 0.117647
K_8 X_COLL_1.L_CORE X_COLL_3.L_CORE 0.058824
K_9 X_COLL_1.L_CORE X_COLL_4.L_CORE 0.117647
K_10 X_COLL_1.L_CORE X_COLL_5.L_CORE 0.083189
K_11 X_COLL_1.L_CORE X_COLL_6.L_CORE 0.052613
K_12 X_COLL_1.L_CORE X_COLL_7.L_CORE 0.058824
K_13 X_COLL_1.L_CORE X_COLL_8.L_CORE 0.052613
K_14 X_COLL_1.L_CORE X_COLL_9.L_CORE 0.041595
K_15 X_COLL_2.L_CORE X_COLL_3.L_CORE 0.117647
K_16 X_COLL_2.L_CORE X_COLL_4.L_CORE 0.083189
K_17 X_COLL_2.L_CORE X_COLL_5.L_CORE 0.117647
K_18 X_COLL_2.L_CORE X_COLL_6.L_CORE 0.083189
K_19 X_COLL_2.L_CORE X_COLL_7.L_CORE 0.052613
K_20 X_COLL_2.L_CORE X_COLL_8.L_CORE 0.058824
K_21 X_COLL_2.L_CORE X_COLL_9.L_CORE 0.052613
K_22 X_COLL_3.L_CORE X_COLL_4.L_CORE 0.052613
K_23 X_COLL_3.L_CORE X_COLL_5.L_CORE 0.083189
K_24 X_COLL_3.L_CORE X_COLL_6.L_CORE 0.117647
K_25 X_COLL_3.L_CORE X_COLL_7.L_CORE 0.041595
K_26 X_COLL_3.L_CORE X_COLL_8.L_CORE 0.052613
K_27 X_COLL_3.L_CORE X_COLL_9.L_CORE 0.058824
K_28 X_COLL_4.L_CORE X_COLL_5.L_CORE 0.117647
K_29 X_COLL_4.L_CORE X_COLL_6.L_CORE 0.058824
K_30 X_COLL_4.L_CORE X_COLL_7.L_CORE 0.117647
K_31 X_COLL_4.L_CORE X_COLL_8.L_CORE 0.083189
K_32 X_COLL_4.L_CORE X_COLL_9.L_CORE 0.052613
K_33 X_COLL_5.L_CORE X_COLL_6.L_CORE 0.117647
K_34 X_COLL_5.L_CORE X_COLL_7.L_CORE 0.083189
K_35 X_COLL_5.L_CORE X_COLL_8.L_CORE 0.117647
K_36 X_COLL_5.L_CORE X_COLL_9.L_CORE 0.083189
K_37 X_COLL_6.L_CORE X_COLL_7.L_CORE 0.052613
K_38 X_COLL_6.L_CORE X_COLL_8.L_CORE 0.083189
K_39 X_COLL_6.L_CORE X_COLL_9.L_CORE 0.117647
K_40 X_COLL_7.L_CORE X_COLL_8.L_CORE 0.117647
K_41 X_COLL_7.L_CORE X_COLL_9.L_CORE 0.058824
K_42 X_COLL_8.L_CORE X_COLL_9.L_CORE 0.117647
* -- Rectification Gradient (Gap Trans-Admittance) --
K_43 X_EMIT_1.L_CORE X_COLL_1.L_CORE 0.011378
K_44 X_EMIT_1.L_CORE X_COLL_2.L_CORE 0.011453
K_45 X_EMIT_1.L_CORE X_COLL_3.L_CORE 0.011420
K_46 X_EMIT_1.L_CORE X_COLL_4.L_CORE 0.011453
K_47 X_EMIT_1.L_CORE X_COLL_5.L_CORE 0.011530
K_48 X_EMIT_1.L_CORE X_COLL_6.L_CORE 0.011497
K_49 X_EMIT_1.L_CORE X_COLL_7.L_CORE 0.011420
K_50 X_EMIT_1.L_CORE X_COLL_8.L_CORE 0.011497
K_51 X_EMIT_1.L_CORE X_COLL_9.L_CORE 0.011464
K_52 X_EMIT_2.L_CORE X_COLL_1.L_CORE 0.011464
K_53 X_EMIT_2.L_CORE X_COLL_2.L_CORE 0.011497
K_54 X_EMIT_2.L_CORE X_COLL_3.L_CORE 0.011420
K_55 X_EMIT_2.L_CORE X_COLL_4.L_CORE 0.011497
K_56 X_EMIT_2.L_CORE X_COLL_5.L_CORE 0.011530
K_57 X_EMIT_2.L_CORE X_COLL_6.L_CORE 0.011453
K_58 X_EMIT_2.L_CORE X_COLL_7.L_CORE 0.011420
K_59 X_EMIT_2.L_CORE X_COLL_8.L_CORE 0.011453
K_60 X_EMIT_2.L_CORE X_COLL_9.L_CORE 0.011378
K_61 X_EMIT_3.L_CORE X_COLL_1.L_CORE 0.011877
K_62 X_EMIT_3.L_CORE X_COLL_2.L_CORE 0.011963
K_63 X_EMIT_3.L_CORE X_COLL_3.L_CORE 0.011926
K_64 X_EMIT_3.L_CORE X_COLL_4.L_CORE 0.011913
K_65 X_EMIT_3.L_CORE X_COLL_5.L_CORE 0.012000
K_66 X_EMIT_3.L_CORE X_COLL_6.L_CORE 0.011963
K_67 X_EMIT_3.L_CORE X_COLL_7.L_CORE 0.011829
K_68 X_EMIT_3.L_CORE X_COLL_8.L_CORE 0.011913
K_69 X_EMIT_3.L_CORE X_COLL_9.L_CORE 0.011877
K_70 X_EMIT_4.L_CORE X_COLL_1.L_CORE 0.011877
K_71 X_EMIT_4.L_CORE X_COLL_2.L_CORE 0.011913
K_72 X_EMIT_4.L_CORE X_COLL_3.L_CORE 0.011829
K_73 X_EMIT_4.L_CORE X_COLL_4.L_CORE 0.011963
K_74 X_EMIT_4.L_CORE X_COLL_5.L_CORE 0.012000
K_75 X_EMIT_4.L_CORE X_COLL_6.L_CORE 0.011913
K_76 X_EMIT_4.L_CORE X_COLL_7.L_CORE 0.011926
K_77 X_EMIT_4.L_CORE X_COLL_8.L_CORE 0.011963
K_78 X_EMIT_4.L_CORE X_COLL_9.L_CORE 0.011877


* -----------------------------------------------------------------
* SIMULATION DIRECTIVES
* -----------------------------------------------------------------
.TRAN 0.1n 50n
* Monitor the inductive momentum coupling across the gap
.PROBE V(NODE_E)

.END
